module top_tb;
    interface aes_if dut_interface;
    
    aes_top DUT(dut_interface);

    

endmodule